-- host.vhd

-- Generated using ACDS version 14.1 190 at 2015.09.10.18:15:58

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity host is
	port (
		atari_d500_byte_export            : in    std_logic_vector(7 downto 0)  := (others => '0'); --         atari_d500_byte.export
		cart_memory_s2_address            : in    std_logic_vector(12 downto 0) := (others => '0'); --          cart_memory_s2.address
		cart_memory_s2_chipselect         : in    std_logic                     := '0';             --                        .chipselect
		cart_memory_s2_clken              : in    std_logic                     := '0';             --                        .clken
		cart_memory_s2_write              : in    std_logic                     := '0';             --                        .write
		cart_memory_s2_readdata           : out   std_logic_vector(7 downto 0);                     --                        .readdata
		cart_memory_s2_writedata          : in    std_logic_vector(7 downto 0)  := (others => '0'); --                        .writedata
		clk_clk                           : in    std_logic                     := '0';             --                     clk.clk
		ext_sram_atari_bus_driven_export  : in    std_logic                     := '0';             --                ext_sram.atari_bus_driven_export
		ext_sram_atari_sram_addr_export   : in    std_logic_vector(19 downto 0) := (others => '0'); --                        .atari_sram_addr_export
		ext_sram_atari_sram_data_export   : out   std_logic_vector(7 downto 0);                     --                        .atari_sram_data_export
		ext_sram_atari_sram_enable_export : in    std_logic                     := '0';             --                        .atari_sram_enable_export
		ext_sram_sram_addr_export         : out   std_logic_vector(19 downto 0);                    --                        .sram_addr_export
		ext_sram_sram_dq_export           : inout std_logic_vector(7 downto 0)  := (others => '0'); --                        .sram_dq_export
		ext_sram_sram_ce_export           : out   std_logic;                                        --                        .sram_ce_export
		ext_sram_sram_oe_n_export         : out   std_logic;                                        --                        .sram_oe_n_export
		ext_sram_sram_we_n_export         : out   std_logic;                                        --                        .sram_we_n_export
		led_external_connection_export    : out   std_logic_vector(4 downto 0);                     -- led_external_connection.export
		reset_reset_n                     : in    std_logic                     := '0';             --                   reset.reset_n
		reset_d500_export                 : out   std_logic;                                        --              reset_d500.export
		sel_cartridge_type_export         : out   std_logic_vector(7 downto 0);                     --      sel_cartridge_type.export
		spi_master_0_cs                   : out   std_logic;                                        --            spi_master_0.cs
		spi_master_0_sclk                 : out   std_logic;                                        --                        .sclk
		spi_master_0_mosi                 : out   std_logic;                                        --                        .mosi
		spi_master_0_miso                 : in    std_logic                     := '0';             --                        .miso
		spi_master_0_cd                   : in    std_logic                     := '0';             --                        .cd
		spi_master_0_wp                   : in    std_logic                     := '0'              --                        .wp
	);
end entity host;

architecture rtl of host is
	component host_atari_d500_byte is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component host_atari_d500_byte;

	component host_cart_memory is
		port (
			address     : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(7 downto 0);                     -- readdata
			writedata   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			address2    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(7 downto 0);                     -- readdata
			writedata2  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X'              -- reset_req
		);
	end component host_cart_memory;

	component host_cpu is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(21 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(21 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component host_cpu;

	component ext_sram_controller is
		port (
			clk               : in    std_logic                     := 'X';             -- clk
			reset             : in    std_logic                     := 'X';             -- reset
			address           : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			chipselect_n      : in    std_logic                     := 'X';             -- chipselect_n
			read_n            : in    std_logic                     := 'X';             -- read_n
			write_n           : in    std_logic                     := 'X';             -- write_n
			writedata         : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			readdata          : out   std_logic_vector(7 downto 0);                     -- readdata
			atari_bus_driven  : in    std_logic                     := 'X';             -- atari_bus_driven_export
			atari_sram_addr   : in    std_logic_vector(19 downto 0) := (others => 'X'); -- atari_sram_addr_export
			atari_sram_data   : out   std_logic_vector(7 downto 0);                     -- atari_sram_data_export
			atari_sram_enable : in    std_logic                     := 'X';             -- atari_sram_enable_export
			sram_addr         : out   std_logic_vector(19 downto 0);                    -- sram_addr_export
			sram_dq           : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- sram_dq_export
			sram_ce           : out   std_logic;                                        -- sram_ce_export
			sram_oe_n         : out   std_logic;                                        -- sram_oe_n_export
			sram_we_n         : out   std_logic                                         -- sram_we_n_export
		);
	end component ext_sram_controller;

	component host_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component host_jtag_uart_0;

	component host_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(4 downto 0)                      -- export
		);
	end component host_led;

	component host_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component host_memory;

	component host_reset_d500 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component host_reset_d500;

	component host_sel_cartridge_type is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component host_sel_cartridge_type;

	component spi_master_if is
		port (
			reset      : in  std_logic                     := 'X';             -- reset
			clk        : in  std_logic                     := 'X';             -- clk
			chipselect : in  std_logic                     := 'X';             -- chipselect
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read       : in  std_logic                     := 'X';             -- read
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			cs         : out std_logic;                                        -- export
			sclk       : out std_logic;                                        -- export
			mosi       : out std_logic;                                        -- export
			miso       : in  std_logic                     := 'X';             -- export
			cd         : in  std_logic                     := 'X';             -- export
			wp         : in  std_logic                     := 'X'              -- export
		);
	end component spi_master_if;

	component host_sysid_2466 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component host_sysid_2466;

	component host_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component host_timer_0;

	component host_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                 : in  std_logic                     := 'X';             -- clk
			cpu_reset_n_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                       : in  std_logic_vector(21 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                   : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                          : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                      : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                         : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                   : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                : in  std_logic_vector(21 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest            : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                   : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			atari_d500_byte_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			atari_d500_byte_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cart_memory_s1_address                        : out std_logic_vector(12 downto 0);                    -- address
			cart_memory_s1_write                          : out std_logic;                                        -- write
			cart_memory_s1_readdata                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			cart_memory_s1_writedata                      : out std_logic_vector(7 downto 0);                     -- writedata
			cart_memory_s1_chipselect                     : out std_logic;                                        -- chipselect
			cart_memory_s1_clken                          : out std_logic;                                        -- clken
			cpu_jtag_debug_module_address                 : out std_logic_vector(8 downto 0);                     -- address
			cpu_jtag_debug_module_write                   : out std_logic;                                        -- write
			cpu_jtag_debug_module_read                    : out std_logic;                                        -- read
			cpu_jtag_debug_module_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_jtag_debug_module_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_jtag_debug_module_byteenable              : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_jtag_debug_module_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			cpu_jtag_debug_module_debugaccess             : out std_logic;                                        -- debugaccess
			ext_sram_controller_0_avalon_slave_address    : out std_logic_vector(19 downto 0);                    -- address
			ext_sram_controller_0_avalon_slave_write      : out std_logic;                                        -- write
			ext_sram_controller_0_avalon_slave_read       : out std_logic;                                        -- read
			ext_sram_controller_0_avalon_slave_readdata   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			ext_sram_controller_0_avalon_slave_writedata  : out std_logic_vector(7 downto 0);                     -- writedata
			ext_sram_controller_0_avalon_slave_chipselect : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address         : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write           : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read            : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect      : out std_logic;                                        -- chipselect
			led_s1_address                                : out std_logic_vector(1 downto 0);                     -- address
			led_s1_write                                  : out std_logic;                                        -- write
			led_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			led_s1_chipselect                             : out std_logic;                                        -- chipselect
			memory_s1_address                             : out std_logic_vector(12 downto 0);                    -- address
			memory_s1_write                               : out std_logic;                                        -- write
			memory_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			memory_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			memory_s1_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			memory_s1_chipselect                          : out std_logic;                                        -- chipselect
			memory_s1_clken                               : out std_logic;                                        -- clken
			reset_d500_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			reset_d500_s1_write                           : out std_logic;                                        -- write
			reset_d500_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			reset_d500_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			reset_d500_s1_chipselect                      : out std_logic;                                        -- chipselect
			sel_cartridge_type_s1_address                 : out std_logic_vector(1 downto 0);                     -- address
			sel_cartridge_type_s1_write                   : out std_logic;                                        -- write
			sel_cartridge_type_s1_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sel_cartridge_type_s1_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			sel_cartridge_type_s1_chipselect              : out std_logic;                                        -- chipselect
			spi_master_0_s1_address                       : out std_logic_vector(2 downto 0);                     -- address
			spi_master_0_s1_write                         : out std_logic;                                        -- write
			spi_master_0_s1_read                          : out std_logic;                                        -- read
			spi_master_0_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			spi_master_0_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			spi_master_0_s1_chipselect                    : out std_logic;                                        -- chipselect
			sysid_2466_control_slave_address              : out std_logic_vector(0 downto 0);                     -- address
			sysid_2466_control_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                            : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                              : out std_logic;                                        -- write
			timer_0_s1_readdata                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                          : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                         : out std_logic                                         -- chipselect
		);
	end component host_mm_interconnect_0;

	component host_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component host_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal cpu_data_master_readdata                                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                               : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                               : std_logic;                     -- cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                                   : std_logic_vector(21 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                                : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                      : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                                     : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                                 : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                        : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                            : std_logic_vector(21 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                               : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect                : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata                  : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest               : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address                   : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                     : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_ext_sram_controller_0_avalon_slave_chipselect           : std_logic;                     -- mm_interconnect_0:ext_sram_controller_0_avalon_slave_chipselect -> mm_interconnect_0_ext_sram_controller_0_avalon_slave_chipselect:in
	signal mm_interconnect_0_ext_sram_controller_0_avalon_slave_readdata             : std_logic_vector(7 downto 0);  -- ext_sram_controller_0:readdata -> mm_interconnect_0:ext_sram_controller_0_avalon_slave_readdata
	signal mm_interconnect_0_ext_sram_controller_0_avalon_slave_address              : std_logic_vector(19 downto 0); -- mm_interconnect_0:ext_sram_controller_0_avalon_slave_address -> ext_sram_controller_0:address
	signal mm_interconnect_0_ext_sram_controller_0_avalon_slave_read                 : std_logic;                     -- mm_interconnect_0:ext_sram_controller_0_avalon_slave_read -> mm_interconnect_0_ext_sram_controller_0_avalon_slave_read:in
	signal mm_interconnect_0_ext_sram_controller_0_avalon_slave_write                : std_logic;                     -- mm_interconnect_0:ext_sram_controller_0_avalon_slave_write -> mm_interconnect_0_ext_sram_controller_0_avalon_slave_write:in
	signal mm_interconnect_0_ext_sram_controller_0_avalon_slave_writedata            : std_logic_vector(7 downto 0);  -- mm_interconnect_0:ext_sram_controller_0_avalon_slave_writedata -> ext_sram_controller_0:writedata
	signal mm_interconnect_0_sysid_2466_control_slave_readdata                       : std_logic_vector(31 downto 0); -- sysid_2466:readdata -> mm_interconnect_0:sysid_2466_control_slave_readdata
	signal mm_interconnect_0_sysid_2466_control_slave_address                        : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_2466_control_slave_address -> sysid_2466:address
	signal mm_interconnect_0_cpu_jtag_debug_module_readdata                          : std_logic_vector(31 downto 0); -- cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	signal mm_interconnect_0_cpu_jtag_debug_module_waitrequest                       : std_logic;                     -- cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	signal mm_interconnect_0_cpu_jtag_debug_module_debugaccess                       : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	signal mm_interconnect_0_cpu_jtag_debug_module_address                           : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	signal mm_interconnect_0_cpu_jtag_debug_module_read                              : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	signal mm_interconnect_0_cpu_jtag_debug_module_byteenable                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	signal mm_interconnect_0_cpu_jtag_debug_module_write                             : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	signal mm_interconnect_0_cpu_jtag_debug_module_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	signal mm_interconnect_0_memory_s1_chipselect                                    : std_logic;                     -- mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	signal mm_interconnect_0_memory_s1_readdata                                      : std_logic_vector(31 downto 0); -- memory:readdata -> mm_interconnect_0:memory_s1_readdata
	signal mm_interconnect_0_memory_s1_address                                       : std_logic_vector(12 downto 0); -- mm_interconnect_0:memory_s1_address -> memory:address
	signal mm_interconnect_0_memory_s1_byteenable                                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	signal mm_interconnect_0_memory_s1_write                                         : std_logic;                     -- mm_interconnect_0:memory_s1_write -> memory:write
	signal mm_interconnect_0_memory_s1_writedata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:memory_s1_writedata -> memory:writedata
	signal mm_interconnect_0_memory_s1_clken                                         : std_logic;                     -- mm_interconnect_0:memory_s1_clken -> memory:clken
	signal mm_interconnect_0_led_s1_chipselect                                       : std_logic;                     -- mm_interconnect_0:led_s1_chipselect -> led:chipselect
	signal mm_interconnect_0_led_s1_readdata                                         : std_logic_vector(31 downto 0); -- led:readdata -> mm_interconnect_0:led_s1_readdata
	signal mm_interconnect_0_led_s1_address                                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_s1_address -> led:address
	signal mm_interconnect_0_led_s1_write                                            : std_logic;                     -- mm_interconnect_0:led_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_writedata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_s1_writedata -> led:writedata
	signal mm_interconnect_0_timer_0_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                                     : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                                      : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                                        : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_cart_memory_s1_chipselect                               : std_logic;                     -- mm_interconnect_0:cart_memory_s1_chipselect -> cart_memory:chipselect
	signal mm_interconnect_0_cart_memory_s1_readdata                                 : std_logic_vector(7 downto 0);  -- cart_memory:readdata -> mm_interconnect_0:cart_memory_s1_readdata
	signal mm_interconnect_0_cart_memory_s1_address                                  : std_logic_vector(12 downto 0); -- mm_interconnect_0:cart_memory_s1_address -> cart_memory:address
	signal mm_interconnect_0_cart_memory_s1_write                                    : std_logic;                     -- mm_interconnect_0:cart_memory_s1_write -> cart_memory:write
	signal mm_interconnect_0_cart_memory_s1_writedata                                : std_logic_vector(7 downto 0);  -- mm_interconnect_0:cart_memory_s1_writedata -> cart_memory:writedata
	signal mm_interconnect_0_cart_memory_s1_clken                                    : std_logic;                     -- mm_interconnect_0:cart_memory_s1_clken -> cart_memory:clken
	signal mm_interconnect_0_sel_cartridge_type_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:sel_cartridge_type_s1_chipselect -> sel_cartridge_type:chipselect
	signal mm_interconnect_0_sel_cartridge_type_s1_readdata                          : std_logic_vector(31 downto 0); -- sel_cartridge_type:readdata -> mm_interconnect_0:sel_cartridge_type_s1_readdata
	signal mm_interconnect_0_sel_cartridge_type_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sel_cartridge_type_s1_address -> sel_cartridge_type:address
	signal mm_interconnect_0_sel_cartridge_type_s1_write                             : std_logic;                     -- mm_interconnect_0:sel_cartridge_type_s1_write -> mm_interconnect_0_sel_cartridge_type_s1_write:in
	signal mm_interconnect_0_sel_cartridge_type_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:sel_cartridge_type_s1_writedata -> sel_cartridge_type:writedata
	signal mm_interconnect_0_spi_master_0_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:spi_master_0_s1_chipselect -> spi_master_0:chipselect
	signal mm_interconnect_0_spi_master_0_s1_readdata                                : std_logic_vector(31 downto 0); -- spi_master_0:readdata -> mm_interconnect_0:spi_master_0_s1_readdata
	signal mm_interconnect_0_spi_master_0_s1_address                                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_master_0_s1_address -> spi_master_0:address
	signal mm_interconnect_0_spi_master_0_s1_read                                    : std_logic;                     -- mm_interconnect_0:spi_master_0_s1_read -> spi_master_0:read
	signal mm_interconnect_0_spi_master_0_s1_write                                   : std_logic;                     -- mm_interconnect_0:spi_master_0_s1_write -> spi_master_0:write
	signal mm_interconnect_0_spi_master_0_s1_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:spi_master_0_s1_writedata -> spi_master_0:writedata
	signal mm_interconnect_0_atari_d500_byte_s1_readdata                             : std_logic_vector(31 downto 0); -- atari_d500_byte:readdata -> mm_interconnect_0:atari_d500_byte_s1_readdata
	signal mm_interconnect_0_atari_d500_byte_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:atari_d500_byte_s1_address -> atari_d500_byte:address
	signal mm_interconnect_0_reset_d500_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:reset_d500_s1_chipselect -> reset_d500:chipselect
	signal mm_interconnect_0_reset_d500_s1_readdata                                  : std_logic_vector(31 downto 0); -- reset_d500:readdata -> mm_interconnect_0:reset_d500_s1_readdata
	signal mm_interconnect_0_reset_d500_s1_address                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:reset_d500_s1_address -> reset_d500:address
	signal mm_interconnect_0_reset_d500_s1_write                                     : std_logic;                     -- mm_interconnect_0:reset_d500_s1_write -> mm_interconnect_0_reset_d500_s1_write:in
	signal mm_interconnect_0_reset_d500_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:reset_d500_s1_writedata -> reset_d500:writedata
	signal irq_mapper_receiver0_irq                                                  : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                  : std_logic;                     -- timer_0:irq -> irq_mapper:receiver1_irq
	signal cpu_d_irq_irq                                                             : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:d_irq
	signal rst_controller_reset_out_reset                                            : std_logic;                     -- rst_controller:reset_out -> [cart_memory:reset, ext_sram_controller_0:reset, irq_mapper:reset, memory:reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, spi_master_0:reset]
	signal rst_controller_reset_out_reset_req                                        : std_logic;                     -- rst_controller:reset_req -> [cart_memory:reset_req, cpu:reset_req, memory:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                                   : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv            : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv           : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_ext_sram_controller_0_avalon_slave_chipselect_ports_inv : std_logic;                     -- mm_interconnect_0_ext_sram_controller_0_avalon_slave_chipselect:inv -> ext_sram_controller_0:chipselect_n
	signal mm_interconnect_0_ext_sram_controller_0_avalon_slave_read_ports_inv       : std_logic;                     -- mm_interconnect_0_ext_sram_controller_0_avalon_slave_read:inv -> ext_sram_controller_0:read_n
	signal mm_interconnect_0_ext_sram_controller_0_avalon_slave_write_ports_inv      : std_logic;                     -- mm_interconnect_0_ext_sram_controller_0_avalon_slave_write:inv -> ext_sram_controller_0:write_n
	signal mm_interconnect_0_led_s1_write_ports_inv                                  : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> led:write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_sel_cartridge_type_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_sel_cartridge_type_s1_write:inv -> sel_cartridge_type:write_n
	signal mm_interconnect_0_reset_d500_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_reset_d500_s1_write:inv -> reset_d500:write_n
	signal rst_controller_reset_out_reset_ports_inv                                  : std_logic;                     -- rst_controller_reset_out_reset:inv -> [atari_d500_byte:reset_n, cpu:reset_n, jtag_uart_0:rst_n, led:reset_n, reset_d500:reset_n, sel_cartridge_type:reset_n, sysid_2466:reset_n, timer_0:reset_n]

begin

	atari_d500_byte : component host_atari_d500_byte
		port map (
			clk      => clk_clk,                                       --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address  => mm_interconnect_0_atari_d500_byte_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_atari_d500_byte_s1_readdata, --                    .readdata
			in_port  => atari_d500_byte_export                         -- external_connection.export
		);

	cart_memory : component host_cart_memory
		port map (
			address     => mm_interconnect_0_cart_memory_s1_address,    --     s1.address
			clken       => mm_interconnect_0_cart_memory_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_cart_memory_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_cart_memory_s1_write,      --       .write
			readdata    => mm_interconnect_0_cart_memory_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_cart_memory_s1_writedata,  --       .writedata
			address2    => cart_memory_s2_address,                      --     s2.address
			chipselect2 => cart_memory_s2_chipselect,                   --       .chipselect
			clken2      => cart_memory_s2_clken,                        --       .clken
			write2      => cart_memory_s2_write,                        --       .write
			readdata2   => cart_memory_s2_readdata,                     --       .readdata
			writedata2  => cart_memory_s2_writedata,                    --       .writedata
			clk         => clk_clk,                                     --   clk1.clk
			reset       => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req           --       .reset_req
		);

	cpu : component host_cpu
		port map (
			clk                                   => clk_clk,                                             --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,            --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                             => cpu_data_master_address,                             --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                          --                          .byteenable
			d_read                                => cpu_data_master_read,                                --                          .read
			d_readdata                            => cpu_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => cpu_data_master_write,                               --                          .write
			d_writedata                           => cpu_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                      --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                         --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => cpu_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_cpu_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_cpu_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_cpu_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_cpu_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_cpu_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_cpu_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_cpu_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_cpu_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                 -- custom_instruction_master.readra
		);

	ext_sram_controller_0 : component ext_sram_controller
		port map (
			clk               => clk_clk,                                                                   --        clock.clk
			reset             => rst_controller_reset_out_reset,                                            --        reset.reset
			address           => mm_interconnect_0_ext_sram_controller_0_avalon_slave_address,              -- avalon_slave.address
			chipselect_n      => mm_interconnect_0_ext_sram_controller_0_avalon_slave_chipselect_ports_inv, --             .chipselect_n
			read_n            => mm_interconnect_0_ext_sram_controller_0_avalon_slave_read_ports_inv,       --             .read_n
			write_n           => mm_interconnect_0_ext_sram_controller_0_avalon_slave_write_ports_inv,      --             .write_n
			writedata         => mm_interconnect_0_ext_sram_controller_0_avalon_slave_writedata,            --             .writedata
			readdata          => mm_interconnect_0_ext_sram_controller_0_avalon_slave_readdata,             --             .readdata
			atari_bus_driven  => ext_sram_atari_bus_driven_export,                                          --      conduit.atari_bus_driven_export
			atari_sram_addr   => ext_sram_atari_sram_addr_export,                                           --             .atari_sram_addr_export
			atari_sram_data   => ext_sram_atari_sram_data_export,                                           --             .atari_sram_data_export
			atari_sram_enable => ext_sram_atari_sram_enable_export,                                         --             .atari_sram_enable_export
			sram_addr         => ext_sram_sram_addr_export,                                                 --             .sram_addr_export
			sram_dq           => ext_sram_sram_dq_export,                                                   --             .sram_dq_export
			sram_ce           => ext_sram_sram_ce_export,                                                   --             .sram_ce_export
			sram_oe_n         => ext_sram_sram_oe_n_export,                                                 --             .sram_oe_n_export
			sram_we_n         => ext_sram_sram_we_n_export                                                  --             .sram_we_n_export
		);

	jtag_uart_0 : component host_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	led : component host_led
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,        --                    .readdata
			out_port   => led_external_connection_export            -- external_connection.export
		);

	memory : component host_memory
		port map (
			clk        => clk_clk,                                --   clk1.clk
			address    => mm_interconnect_0_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,         -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req      --       .reset_req
		);

	reset_d500 : component host_reset_d500
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_reset_d500_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_reset_d500_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_reset_d500_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_reset_d500_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_reset_d500_s1_readdata,        --                    .readdata
			out_port   => reset_d500_export                                -- external_connection.export
		);

	sel_cartridge_type : component host_sel_cartridge_type
		port map (
			clk        => clk_clk,                                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                --               reset.reset_n
			address    => mm_interconnect_0_sel_cartridge_type_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_sel_cartridge_type_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_sel_cartridge_type_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_sel_cartridge_type_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_sel_cartridge_type_s1_readdata,        --                    .readdata
			out_port   => sel_cartridge_type_export                                -- external_connection.export
		);

	spi_master_0 : component spi_master_if
		port map (
			reset      => rst_controller_reset_out_reset,               --    reset.reset
			clk        => clk_clk,                                      --      clk.clk
			chipselect => mm_interconnect_0_spi_master_0_s1_chipselect, --       s1.chipselect
			address    => mm_interconnect_0_spi_master_0_s1_address,    --         .address
			write      => mm_interconnect_0_spi_master_0_s1_write,      --         .write
			writedata  => mm_interconnect_0_spi_master_0_s1_writedata,  --         .writedata
			read       => mm_interconnect_0_spi_master_0_s1_read,       --         .read
			readdata   => mm_interconnect_0_spi_master_0_s1_readdata,   --         .readdata
			cs         => spi_master_0_cs,                              -- external.export
			sclk       => spi_master_0_sclk,                            --         .export
			mosi       => spi_master_0_mosi,                            --         .export
			miso       => spi_master_0_miso,                            --         .export
			cd         => spi_master_0_cd,                              --         .export
			wp         => spi_master_0_wp                               --         .export
		);

	sysid_2466 : component host_sysid_2466
		port map (
			clock    => clk_clk,                                               --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,              --         reset.reset_n
			readdata => mm_interconnect_0_sysid_2466_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_2466_control_slave_address(0)  --              .address
		);

	timer_0 : component host_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	mm_interconnect_0 : component host_mm_interconnect_0
		port map (
			clk_0_clk_clk                                 => clk_clk,                                                         --                          clk_0_clk.clk
			cpu_reset_n_reset_bridge_in_reset_reset       => rst_controller_reset_out_reset,                                  --  cpu_reset_n_reset_bridge_in_reset.reset
			cpu_data_master_address                       => cpu_data_master_address,                                         --                    cpu_data_master.address
			cpu_data_master_waitrequest                   => cpu_data_master_waitrequest,                                     --                                   .waitrequest
			cpu_data_master_byteenable                    => cpu_data_master_byteenable,                                      --                                   .byteenable
			cpu_data_master_read                          => cpu_data_master_read,                                            --                                   .read
			cpu_data_master_readdata                      => cpu_data_master_readdata,                                        --                                   .readdata
			cpu_data_master_write                         => cpu_data_master_write,                                           --                                   .write
			cpu_data_master_writedata                     => cpu_data_master_writedata,                                       --                                   .writedata
			cpu_data_master_debugaccess                   => cpu_data_master_debugaccess,                                     --                                   .debugaccess
			cpu_instruction_master_address                => cpu_instruction_master_address,                                  --             cpu_instruction_master.address
			cpu_instruction_master_waitrequest            => cpu_instruction_master_waitrequest,                              --                                   .waitrequest
			cpu_instruction_master_read                   => cpu_instruction_master_read,                                     --                                   .read
			cpu_instruction_master_readdata               => cpu_instruction_master_readdata,                                 --                                   .readdata
			atari_d500_byte_s1_address                    => mm_interconnect_0_atari_d500_byte_s1_address,                    --                 atari_d500_byte_s1.address
			atari_d500_byte_s1_readdata                   => mm_interconnect_0_atari_d500_byte_s1_readdata,                   --                                   .readdata
			cart_memory_s1_address                        => mm_interconnect_0_cart_memory_s1_address,                        --                     cart_memory_s1.address
			cart_memory_s1_write                          => mm_interconnect_0_cart_memory_s1_write,                          --                                   .write
			cart_memory_s1_readdata                       => mm_interconnect_0_cart_memory_s1_readdata,                       --                                   .readdata
			cart_memory_s1_writedata                      => mm_interconnect_0_cart_memory_s1_writedata,                      --                                   .writedata
			cart_memory_s1_chipselect                     => mm_interconnect_0_cart_memory_s1_chipselect,                     --                                   .chipselect
			cart_memory_s1_clken                          => mm_interconnect_0_cart_memory_s1_clken,                          --                                   .clken
			cpu_jtag_debug_module_address                 => mm_interconnect_0_cpu_jtag_debug_module_address,                 --              cpu_jtag_debug_module.address
			cpu_jtag_debug_module_write                   => mm_interconnect_0_cpu_jtag_debug_module_write,                   --                                   .write
			cpu_jtag_debug_module_read                    => mm_interconnect_0_cpu_jtag_debug_module_read,                    --                                   .read
			cpu_jtag_debug_module_readdata                => mm_interconnect_0_cpu_jtag_debug_module_readdata,                --                                   .readdata
			cpu_jtag_debug_module_writedata               => mm_interconnect_0_cpu_jtag_debug_module_writedata,               --                                   .writedata
			cpu_jtag_debug_module_byteenable              => mm_interconnect_0_cpu_jtag_debug_module_byteenable,              --                                   .byteenable
			cpu_jtag_debug_module_waitrequest             => mm_interconnect_0_cpu_jtag_debug_module_waitrequest,             --                                   .waitrequest
			cpu_jtag_debug_module_debugaccess             => mm_interconnect_0_cpu_jtag_debug_module_debugaccess,             --                                   .debugaccess
			ext_sram_controller_0_avalon_slave_address    => mm_interconnect_0_ext_sram_controller_0_avalon_slave_address,    -- ext_sram_controller_0_avalon_slave.address
			ext_sram_controller_0_avalon_slave_write      => mm_interconnect_0_ext_sram_controller_0_avalon_slave_write,      --                                   .write
			ext_sram_controller_0_avalon_slave_read       => mm_interconnect_0_ext_sram_controller_0_avalon_slave_read,       --                                   .read
			ext_sram_controller_0_avalon_slave_readdata   => mm_interconnect_0_ext_sram_controller_0_avalon_slave_readdata,   --                                   .readdata
			ext_sram_controller_0_avalon_slave_writedata  => mm_interconnect_0_ext_sram_controller_0_avalon_slave_writedata,  --                                   .writedata
			ext_sram_controller_0_avalon_slave_chipselect => mm_interconnect_0_ext_sram_controller_0_avalon_slave_chipselect, --                                   .chipselect
			jtag_uart_0_avalon_jtag_slave_address         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,         --      jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,           --                                   .write
			jtag_uart_0_avalon_jtag_slave_read            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,            --                                   .read
			jtag_uart_0_avalon_jtag_slave_readdata        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                                   .readdata
			jtag_uart_0_avalon_jtag_slave_writedata       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                                   .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                                   .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      --                                   .chipselect
			led_s1_address                                => mm_interconnect_0_led_s1_address,                                --                             led_s1.address
			led_s1_write                                  => mm_interconnect_0_led_s1_write,                                  --                                   .write
			led_s1_readdata                               => mm_interconnect_0_led_s1_readdata,                               --                                   .readdata
			led_s1_writedata                              => mm_interconnect_0_led_s1_writedata,                              --                                   .writedata
			led_s1_chipselect                             => mm_interconnect_0_led_s1_chipselect,                             --                                   .chipselect
			memory_s1_address                             => mm_interconnect_0_memory_s1_address,                             --                          memory_s1.address
			memory_s1_write                               => mm_interconnect_0_memory_s1_write,                               --                                   .write
			memory_s1_readdata                            => mm_interconnect_0_memory_s1_readdata,                            --                                   .readdata
			memory_s1_writedata                           => mm_interconnect_0_memory_s1_writedata,                           --                                   .writedata
			memory_s1_byteenable                          => mm_interconnect_0_memory_s1_byteenable,                          --                                   .byteenable
			memory_s1_chipselect                          => mm_interconnect_0_memory_s1_chipselect,                          --                                   .chipselect
			memory_s1_clken                               => mm_interconnect_0_memory_s1_clken,                               --                                   .clken
			reset_d500_s1_address                         => mm_interconnect_0_reset_d500_s1_address,                         --                      reset_d500_s1.address
			reset_d500_s1_write                           => mm_interconnect_0_reset_d500_s1_write,                           --                                   .write
			reset_d500_s1_readdata                        => mm_interconnect_0_reset_d500_s1_readdata,                        --                                   .readdata
			reset_d500_s1_writedata                       => mm_interconnect_0_reset_d500_s1_writedata,                       --                                   .writedata
			reset_d500_s1_chipselect                      => mm_interconnect_0_reset_d500_s1_chipselect,                      --                                   .chipselect
			sel_cartridge_type_s1_address                 => mm_interconnect_0_sel_cartridge_type_s1_address,                 --              sel_cartridge_type_s1.address
			sel_cartridge_type_s1_write                   => mm_interconnect_0_sel_cartridge_type_s1_write,                   --                                   .write
			sel_cartridge_type_s1_readdata                => mm_interconnect_0_sel_cartridge_type_s1_readdata,                --                                   .readdata
			sel_cartridge_type_s1_writedata               => mm_interconnect_0_sel_cartridge_type_s1_writedata,               --                                   .writedata
			sel_cartridge_type_s1_chipselect              => mm_interconnect_0_sel_cartridge_type_s1_chipselect,              --                                   .chipselect
			spi_master_0_s1_address                       => mm_interconnect_0_spi_master_0_s1_address,                       --                    spi_master_0_s1.address
			spi_master_0_s1_write                         => mm_interconnect_0_spi_master_0_s1_write,                         --                                   .write
			spi_master_0_s1_read                          => mm_interconnect_0_spi_master_0_s1_read,                          --                                   .read
			spi_master_0_s1_readdata                      => mm_interconnect_0_spi_master_0_s1_readdata,                      --                                   .readdata
			spi_master_0_s1_writedata                     => mm_interconnect_0_spi_master_0_s1_writedata,                     --                                   .writedata
			spi_master_0_s1_chipselect                    => mm_interconnect_0_spi_master_0_s1_chipselect,                    --                                   .chipselect
			sysid_2466_control_slave_address              => mm_interconnect_0_sysid_2466_control_slave_address,              --           sysid_2466_control_slave.address
			sysid_2466_control_slave_readdata             => mm_interconnect_0_sysid_2466_control_slave_readdata,             --                                   .readdata
			timer_0_s1_address                            => mm_interconnect_0_timer_0_s1_address,                            --                         timer_0_s1.address
			timer_0_s1_write                              => mm_interconnect_0_timer_0_s1_write,                              --                                   .write
			timer_0_s1_readdata                           => mm_interconnect_0_timer_0_s1_readdata,                           --                                   .readdata
			timer_0_s1_writedata                          => mm_interconnect_0_timer_0_s1_writedata,                          --                                   .writedata
			timer_0_s1_chipselect                         => mm_interconnect_0_timer_0_s1_chipselect                          --                                   .chipselect
		);

	irq_mapper : component host_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_d_irq_irq                   --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_ext_sram_controller_0_avalon_slave_chipselect_ports_inv <= not mm_interconnect_0_ext_sram_controller_0_avalon_slave_chipselect;

	mm_interconnect_0_ext_sram_controller_0_avalon_slave_read_ports_inv <= not mm_interconnect_0_ext_sram_controller_0_avalon_slave_read;

	mm_interconnect_0_ext_sram_controller_0_avalon_slave_write_ports_inv <= not mm_interconnect_0_ext_sram_controller_0_avalon_slave_write;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_sel_cartridge_type_s1_write_ports_inv <= not mm_interconnect_0_sel_cartridge_type_s1_write;

	mm_interconnect_0_reset_d500_s1_write_ports_inv <= not mm_interconnect_0_reset_d500_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of host
